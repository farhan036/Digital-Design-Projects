

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO SYS_TOP 
  PIN SI[3] 
    ANTENNAPARTIALMETALAREA 0.228 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.09668 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.368 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.96248 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32756 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 23.533 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 113.386 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 625.453 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 3022.22 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 4.74109 LAYER VIA56 ;
  END SI[3]
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 0.816 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.92496 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.268 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48148 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 32.33 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 155.7 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 645.791 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 3120.04 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 4.06379 LAYER VIA56 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 0.438 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.10678 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.286 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1881 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.117 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.2352 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 4.523 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.948 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 136.992 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 672.717 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.38649 LAYER VIA56 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 2.005 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.64405 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.359 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1592 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 90.5375 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 442.054 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA34 ;
  END SI[0]
  PIN SO[3] 
    ANTENNADIFFAREA 0.537 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 6.155 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.6056 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 48.5336 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 231.881 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.53405 LAYER VIA34 ;
  END SO[3]
  PIN SO[2] 
    ANTENNAPARTIALMETALAREA 2.789 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.4151 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 32.412 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 156.094 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 181.186 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 873.633 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.90476 LAYER VIA56 ;
  END SO[2]
  PIN SO[1] 
    ANTENNAPARTIALMETALAREA 0.487 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.34247 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.25 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3949 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 29.214 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 140.712 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8216 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 53.8197 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 257.832 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.878773 LAYER VIA56 ;
  END SO[1]
  PIN SO[0] 
    ANTENNAPARTIALMETALAREA 2.179 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.481 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.386 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 40.5291 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 124.069 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 602.394 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.90126 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 29.36 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 141.414 LAYER METAL5 ;
    ANTENNAGATEAREA 0.2171 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 259.306 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1253.77 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 4.17746 LAYER VIA56 ;
  END SO[0]
  PIN SE 
    ANTENNAPARTIALMETALAREA 1.995 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.59595 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.099 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.9086 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1755 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 27.7869 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 135.072 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.411396 LAYER VIA34 ;
  END SE
  PIN scan_clk 
    ANTENNAPARTIALMETALAREA 0.255 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.22655 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.878 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.41558 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.206 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.99326 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 0.735144 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 3.68179 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END scan_clk
  PIN scan_rst 
    ANTENNAPARTIALMETALAREA 1.353 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.50793 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.751 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.80471 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 11.01 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 53.1505 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 305.872 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1478.61 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 4.06379 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 13.151 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 63.4487 LAYER METAL5 ;
    ANTENNAGATEAREA 0.1599 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 388.118 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1875.41 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 4.74109 LAYER VIA56 ;
  END scan_rst
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 0.551 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.65031 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.525 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1477 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 44.6774 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 218.312 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.828932 LAYER VIA34 ;
  END test_mode
  PIN REF_CLK 
    ANTENNAPARTIALMETALAREA 0.619 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.97739 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.698 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.35978 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 0.689434 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 3.39911 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END REF_CLK
  PIN UART_CLK 
    ANTENNAPARTIALMETALAREA 0.241 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.15921 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.206 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.99326 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.62674 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 0.60128 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 3.0379 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END UART_CLK
  PIN RST_N 
    ANTENNAPARTIALMETALAREA 0.893 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.29533 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.25 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3949 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.928 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 43.1361 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 326.979 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1580.13 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA45 ;
  END RST_N
  PIN UART_RX_IN 
    ANTENNAPARTIALMETALAREA 1.586 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.62866 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 19.866 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 95.7479 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5057 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 50.4213 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 242.728 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 1.42675 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 9.689 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 46.7965 LAYER METAL5 ;
    ANTENNAGATEAREA 0.7111 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 64.0467 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 308.536 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.42675 LAYER VIA56 ;
  END UART_RX_IN
  PIN UART_TX_O 
    ANTENNAPARTIALMETALAREA 11.444 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.0456 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.213 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8369 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 1.529 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 9.206 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 44.4733 LAYER METAL5 ;
  END UART_TX_O
  PIN parity_error 
    ANTENNAPARTIALMETALAREA 8.638 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.5488 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 11.971 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 57.7729 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 26.344 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 126.907 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3185 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 193.247 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 935.497 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.83987 LAYER VIA56 ;
  END parity_error
  PIN framing_error 
    ANTENNADIFFAREA 0.524 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.807 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.88167 LAYER METAL3 ;
  END framing_error
END SYS_TOP

END LIBRARY
