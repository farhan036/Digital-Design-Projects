module FSM (
    input wire        CLK,
    input wire        RST,          // Asynchronous Active Low Reset
    input wire        RX_IN,        // Serial input line
    input wire        PAR_EN,       // Parity enable
    input wire  [3:0] bit_cnt,      // Bit counter
    input wire  [4:0] edge_cnt,     // Edge counter 
    input  wire [5:0] Prescale,     // Sampling rate: 8, 16, 32
    input wire        par_err,      // Parity error flag
    input wire        strt_glitch,  // Start glitch detected
    input wire        stp_err,      // Stop bit error flag
    output reg        par_chk_en,   // Enable parity check
    output reg        strt_chk_en,  // Enable start check
    output reg        stp_chk_en,   // Enable stop check
    output reg        enable,       // Enable edge/bit counter
    output reg        dat_samp_en,  // Enable data sampling
    output reg        deser_en,     // Enable deserializer
    output reg        data_valid    // Data valid pulse (end of frame)
);

    // Gray-coded State Encoding (3-bit)
    typedef enum logic [2:0] {
        IDLE   = 3'b000,
        START  = 3'b001,
        SEND   = 3'b011,
        PARITY = 3'b010,
        STOP   = 3'b110,
        FINAL  = 3'b111
    } state;

    state current_state, next_state;

    //==================================================================
    // Sequential state update
    //==================================================================
    always @(posedge CLK or negedge RST) begin
        if (!RST)
            current_state <= IDLE;
        else
            current_state <= next_state;
    end

    //==================================================================
    // Combinational next-state logic & output control
    //==================================================================
    always @(*) begin
        // Default values
        par_chk_en  = 0;
        strt_chk_en = 0;
        stp_chk_en  = 0;
        enable      = 0;
        dat_samp_en = 0;
        deser_en    = 0;
        data_valid  = 0;

        case (current_state)
            IDLE: begin     // IDLE: Wait for start bit (RX_IN = 0)
                if (RX_IN)
                begin
                    next_state = IDLE;
                end
                else
                    next_state = START;
            end

            START: begin       // START: Sample and validate start bit
                dat_samp_en = 1;    // Enable sampling
                strt_chk_en = 1;    // Enable start check
                enable      = 1;    // Enable edge/bit counter
                if (edge_cnt == Prescale-1 ) 
                begin
                    if (strt_glitch)
                        next_state = IDLE;  // Invalid start bit
                    else
                        next_state = SEND;  // Valid start → receive data
                    end
                else 
                begin
                        next_state = START;
                end
            end

            // SEND: Receive 8 data bits
            SEND: begin
                deser_en    = 1;    // Enable deserializer
                dat_samp_en = 1;    // Enable sampling
                enable      = 1;    // Enable edge/bit counter
                if (bit_cnt == 4'd9) begin
                    if (PAR_EN)
                        next_state = PARITY;    // Go check parity
                    else
                        next_state = STOP;      // Skip to stop bit
                end
                else
                    next_state = SEND;
            end

            // PARITY: Check parity bit (if enabled)
            PARITY: begin
                par_chk_en = 1;     // Enable parity check
                enable     = 1;     // Enable sampling
                dat_samp_en = 1;    // Enable edge/bit counter
                if (bit_cnt == 4'd10)
                begin
                    if(par_err == 1)
                    next_state = IDLE;      // Parity failed → IDLE
                    else
                    next_state = STOP;      // Parity OK → check stop
                end
                else
                    next_state = PARITY;
                
            end

            // STOP: Check stop bit
            STOP: begin
 		  stp_chk_en = 1;     // Enable stop check
                enable     = 1;     // Enable sampling
                dat_samp_en = 1;    // Enable edge/bit counter
                if (PAR_EN) 
                begin
                    if (bit_cnt == 4'd11)
                    begin
                        if(stp_err == 1)
                        next_state = IDLE;      // Stop error → IDLE
                        else
                        next_state = FINAL;     // Stop OK → FINAL
                    end
                    else
                        next_state = STOP;
                end
                else
                begin
                    if (bit_cnt == 4'd10)
                    begin
                        if(stp_err == 1)
                        next_state = IDLE;
                        else
                        next_state = FINAL;
                    end
                else
                        next_state = STOP;
                end
                
            end

            // FINAL: Frame complete  output valid data
            FINAL: begin
                    
                     data_valid = 1;     // Assert valid if no errors
                    if (RX_IN)
                        next_state = IDLE;      // Wait for next frame
                    else
                        next_state = START;     // Immediately start new frame
                
                
                
            end

            default: next_state = IDLE;
        endcase
    end

endmodule
