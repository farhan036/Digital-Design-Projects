module ClkDiv (
    input  wire       I_ref_clk,        // Reference input clock
    input  wire       I_rst_n,          // Active-low asynchronous reset
    input  wire       I_clk_en,         // Clock divider enable
    input  wire [7:0] I_div_ratio,      // Division ratio (must be > 1 for division)
    output wire        o_div_clk        // Divided clock output
);

    // Internal signals
    wire odd;                   // Division ratio odd/even indicator
    wire [7:0] half_toggle;     // Half-period for even divide
    wire [7:0] half_toggle_p;   // Adjusted half-period for odd divide
    reg  [7:0] counter;         // Counter for clock division
    reg        flag;            // Flag to alternate short/long halves in odd divide
    reg div_clk    ;            // Internal divided clock


    assign odd           = I_div_ratio[0];              // Detect if divide ratio is odd
    assign half_toggle   = (I_div_ratio >> 1) - 1;      // For even divide: toggle at half ratio ,i decrement 1 because counter from 0
    assign half_toggle_p = half_toggle + 1;              // For odd divide: alternate between half_toggle and half_toggle + 1

    // Clock divider logic
    always @(posedge I_ref_clk or negedge I_rst_n) begin
        if (!I_rst_n) 
        begin
            // async reset
            div_clk <= 1'b0;
            counter   <= 8'd0;
            flag      <= 1'b0;
        end 
        else if (I_clk_en && (I_div_ratio > 1)) 
        begin
            // enabled and valid ratio
            if (!odd && (counter >= half_toggle)) 
            begin
                // even divide
                div_clk <= ~div_clk;
                counter   <= 8'd0;
            end
            else if (odd && ((counter >= half_toggle  && !flag) ||(counter >= half_toggle_p &&  flag))) 
            begin
                // odd divide (alternate short/long halves)
                div_clk <= ~div_clk;        // Toggle output
                flag      <= ~flag;         // Alternate flag
                counter   <= 8'd0;          // Reset counter
            end
            else 
            begin
                counter <= counter + 1'd1; // Keep counting
            end
        end 
        else 
        begin
            // disabled → force low
            div_clk   <= 'd0;
            counter   <= 8'd0;
            flag      <= 1'b0;
        end
    end
    // Output selection:
    //   - If reset asserted → force low
    //   - If enabled and ratio > 1 → divided clock
    //   - Else → pass reference clock  
   assign o_div_clk = (!I_rst_n) ? I_ref_clk   : ((I_clk_en && (I_div_ratio > 1))) ? div_clk  :  I_ref_clk  ;   
            


endmodule